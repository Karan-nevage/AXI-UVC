//=============================================================================================
// File: axi_sqr.sv
// Description: Defines the UVM sequencer typedef for AXI transactions.
//=============================================================================================

typedef uvm_sequencer#(axi_tx) axi_sqr;
//=============================================================================================
